candle
    input age "Введите ваш возраст: "
    if age >= 18
        print "Доступ разрешен"
    else
        print "Доступ запрещен"
    end
end

[
    Keyword("candle"),
    InstrEnd,
    Atom("input"),
    Atom("age"),
    Quote,
    Atom("Введите"),
    Atom("ваш"),
    Atom("возраст"),
    Atom(":"),
    Quote,
    InstrEnd,
    Keyword("if"),
    Atom("age"),
    Op(
        [
            '>',
        ],
    ),
    Op(
        [
            '=',
        ],
    ),
    Atom(
        [
            '1',
            '8',
        ],
    ),
    InstrEnd,
    Atom(
        [
            'p',
            'r',
            'i',
            'n',
            't',
        ],
    ),
    Quote,
    Atom(
        [
            'Д',
            'о',
            'с',
            'т',
            'у',
            'п',
        ],
    ),
    Atom(
        [
            'р',
            'а',
            'з',
            'р',
            'е',
            'ш',
            'е',
            'н',
        ],
    ),
    Quote,
    InstrEnd,
    Keyword(
        [
            'e',
            'l',
            's',
            'e',
        ],
    ),
    InstrEnd,
    Atom(
        [
            'p',
            'r',
            'i',
            'n',
            't',
        ],
    ),
    Quote,
    Atom(
        [
            'Д',
            'о',
            'с',
            'т',
            'у',
            'п',
        ],
    ),
    Atom(
        [
            'з',
            'а',
            'п',
            'р',
            'е',
            'щ',
            'е',
            'н',
        ],
    ),
    Quote,
    InstrEnd,
    Keyword(
        [
            'e',
            'n',
            'd',
        ],
    ),
    InstrEnd,
    Keyword(
        [
            'e',
            'n',
            'd',
        ],
    ),
    InstrEnd,
]]]Y&*(EHIU(g8yebu987ehiuEHD(*&#RHJ*()#WUR*()#RJ)*RJ$POKopfl=pdl}POEFKJOIFJWIOweh