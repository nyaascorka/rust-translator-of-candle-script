candle
    0nh
endд