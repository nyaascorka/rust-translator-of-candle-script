candle
end